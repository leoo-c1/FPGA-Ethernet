import eth_types_pkg::*

module eth_parser #(
    parameter FPGA_MAC = 48'h00_1A_2B_3C_4D_5E, // FPGA's MAC address (theoretical)
    parameter FPGA_IP = 32'hC0_00_02_92,        // FPGA's IP address (theoretical)
    parameter FPGA_PORT = 16'd5005              // FPGA's UDP port (theoretical)
    ) (
    input logic clk,                    // 50MHz LAN8720 clock
    input logic resetn,                 // Reset button (active low)

    input logic [7:0] received_byte,    // The byte of data we have received from the LAN8720
    input logic byte_valid,             // Pulses for one clock cycle on valid byte

    output logic data,                  // The payload data
    output logic data_valid,            // Whether we are currently sending payload data
    output logic data_last              // Pulses on the last byte of our payload data
    );

    frame_header frame_header_content;  // Each component of the ethernet frame header
    ip_header ip_header_content;        // Each component of the IP packet header
    udp_header udp_header_content;      // Each component of the UDP datagram header

    eth_states state;                   // The current ethernet state we are in

    logic [16:0] ip_checksum_calc;      // The calculated checksum of the IP header
    logic [31:0] ip_checksum_acc;       // 32 bits to handle overflow carries
    logic [15:0] current_word;          // Temporary holder for the 16-bit word

    logic [15:0] byte_counter = 0;      // Counts the number of bytes we have received

    always_ff @ (posedge clk or negedge resetn) begin
        if (!resetn) begin
            state <= IDLE;
            data <= 8'b0;
            data_valid <= 1'b0;
            data_last <= 1'b0;
            byte_counter <= 0;
        end else begin
            if (state == IDLE) begin
                data_valid <= 1'b0;
                data_last <= 1'b0;
                byte_counter <= 0;
                if (byte_valid) begin
                    // If we just received the SFD
                    if (received_byte == 8'hD5)
                        state <= ETH_HEADER;        // Get ready to start reading the frame header
                    else
                        state <= IDLE;
                end else
                    state <= IDLE;
            end else if (state == ETH_HEADER) begin
                // Assign bytes based on the current byte counter
                if (byte_valid) begin
                    if (byte_counter < 6)
                        frame_header_content.dest_mac[byte_counter] <= received_byte;
                    else if (byte_counter < 12)
                        frame_header_content.src_mac[byte_counter-6] <= received_byte;
                    else if (byte_counter < 14)
                        frame_header_content.ethertype[byte_counter-12] <= received_byte;

                    if (byte_counter < 13)
                        byte_counter <= byte_counter + 1;
                    else begin
                        byte_counter <= 0;
                        // Make sure the destination mac is ours and ethertype is 0x0800 (IPv4)
                        if (({>>{frame_header_content.dest_mac}} == FPGA_MAC)
                            & ({frame_header_content.ethertype[0], received_byte} == 16'h0800))
                            state <= IP_HEADER;
                    end
                end

            end else (if state == IP_HEADER) begin
                // Assign bytes based on the current byte counter
                case (byte_counter)
                    0: begin
                        ip_header_content.version <= received_byte[7:4];
                        ip_header_content.header_len <= received_byte[3:0];
                    end

                    1: begin
                        ip_header_content.dscp <= received_byte[7:2];
                        ip_header_content.ecn <= received_byte[1:0];
                    end

                    2: ip_header_content.total_len[0] <= received_byte;
                    3: ip_header_content.total_len[1] <= received_byte;

                    4: ip_header_content.identification[0] <= received_byte;
                    5: ip_header_content.identification[1] <= received_byte;

                    6: begin
                        ip_header_content.flags <= received_byte[7:5];
                        ip_header_content.frag_offset[12:8] <= received_byte[4:0];
                    end
                    7: ip_header_content.frag_offset[7:0] <= received_byte;

                    8: ip_header_content.ttl <= received_byte;

                    9: ip_header_content.protocol <= received_byte;

                    10: ip_header_content.header_csum[0] <= received_byte;
                    11: ip_header_content.header_csum[1] <= received_byte;

                    12: ip_header_content.src_ip[0] <= received_byte;
                    13: ip_header_content.src_ip[1] <= received_byte;
                    14: ip_header_content.src_ip[2] <= received_byte;
                    15: ip_header_content.src_ip[3] <= received_byte;

                    16: ip_header_content.dest_ip[0] <= received_byte;
                    17: ip_header_content.dest_ip[1] <= received_byte;
                    18: ip_header_content.dest_ip[2] <= received_byte;
                    19: ip_header_content.dest_ip[3] <= received_byte;
                endcase

                if (byte_counter[0] == 1'b0) begin
                    // If the current byte is even, it is the MSByte of the 16-bit word
                    current_word[15:8] <= received_byte;
                end 
                else begin
                    // The current byte is odd, so it is the LSByte of the 16-bit word
                    current_word[7:0] <= received_byte;     // Complete the word
                    ip_checksum_acc <= ip_checksum_acc + {current_word[15:8], received_byte};
                end

                if (byte_counter < 19)
                    byte_counter <= byte_counter + 1;
                else begin
                    byte_counter <= 0;

                    // Check if dest_ip matches FPGA's IP
                    if ({ip_header_content.dest_ip[0:2], received_byte} == FPGA_IP)
                        state <= IP_CHECK;
                    else
                        state <= IDLE;
                end
            end else if (state == IP_CHECK) begin
                // Add the carry-over in the checksum to the bottom 16 bits
                ip_checksum_calc <= ip_checksum_acc[31:16] + ip_checksum_acc[15:0];
                // Check if there is still 1 bit of carry-over left over
                if (ip_checksum_calc[16])
                    ip_checksum_calc <= ~(ip_checksum_calc[15:0] + 1'b1);

                // Check if checksum is the valid 0x0000
                if (ip_checksum_calc == 16'h0000)
                    state <= UDP_HEADER;
                else
                    state <= IDLE;

            end else if (state == UDP_HEADER) begin

            end else (if state == PAYLOAD) begin

            end else if (state == FCS) begin

            end else if (state == DONE) begin

            end else begin
                state <= IDLE;
            end
        end
    end

endmodule